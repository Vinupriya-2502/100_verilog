module arithmetic (input a,b,output c);
assign c=a+b;
assign c=a-b;
assign c=a*b;
assign c=a/b;
endmodule
